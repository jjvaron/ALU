library verilog;
use verilog.vl_types.all;
entity multiplicador_vlg_check_tst is
    port(
        product_out     : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end multiplicador_vlg_check_tst;
